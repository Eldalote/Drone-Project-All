library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

entity IMU_compound_filter is
    port (
        clk: in  std_logic;
        rst: in  std_logic
    );
end entity;

architecture rtl of IMU_compound_filter is
begin
end architecture;